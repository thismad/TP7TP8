architecture rtl of collision is

 
  constant x_bat_right : std_logic_vector := "000000000001";  -- pos x of the bat with a -1
  constant x_bat_left  : std_logic_vector := "000000000100"; 
  constant c_compared : std_logic_vector(8 downto 0) := (others => '0');
  signal   s_next_y    : std_logic_vector (8 downto 0);
signal s_and : std_logic_vector (8 downto 0);

begin

  compare : process (x_pos, y_dir)
begin
    if (x_pos = x_bat_right) then
      if (x_dir = '0' and y_dir = '0') then    --bas a gauche
        s_next_y <= y_pos(7 downto 0) & '0';
      elsif(x_dir = '0' and y_dir = '1') then  -- haut gauche
        s_next_y <= '0' & y_pos(8 downto 1);
      end if;
    elsif (x_pos = x_bat_left) then
      if (x_dir = '1' and y_dir = '0') then     --droite haut
        s_next_y <= y_pos(7 downto 0) & '0';
      elsif (x_dir = '1' and y_dir = '1') then  --droite bas
        s_next_y <= '0' & y_pos(8 downto 1);
      end if;
    end if;
  end process;


  tryout : process (x_pos, y_pos, s_and)
  begin
    if(s_and /= c_compared and (x_bat_left = x_pos or x_bat_right = x_pos)) then
      change <= '1';
    else
      change <= '0';
    end if;
  end process;

s_and <= s_next_y and bat_pos;

end architecture rtl;
