architecture rtl of collision is
begin

end architecture rtl;

